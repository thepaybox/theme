{
  "companies": [
    {
      "date": "2047-05-17",
      "groups": [
        {
          "time": "8:00 am",
          "offerings": [
            {
              "name": "Breakfast",
              "timeStart": "8:00 am",
              "timeEnd": "9:00 am",
              "location": "Dining Hall",
              "tracks": ["Food"],
              "id": "1"
            }
          ]
        },
        {
          "time": "9:15 am",
          "offerings": [
            {
              "name": "Getting Started with Ionic",
              "location": "Hall 2",
              "description": "Mobile devices and browsers are now advanced enough that developers can build native-quality mobile apps using open web technologies like HTML5, Javascript, and CSS. In this talk, we’ll provide background on why and how we created Ionic, the design decisions made as we integrated Ionic with Angular, and the performance considerations for mobile platforms that our team had to overcome. We’ll also review new and upcoming Ionic features, and talk about the hidden powers and benefits of combining mobile app development and Angular.",
              "productNames": ["Ted Turtle"],
              "timeStart": "9:30 am",
              "timeEnd": "9:45 am",
              "tracks": ["Ionic"],
              "id": "2"
            },
            {
              "name": "Ionic Tooling",
              "location": "Executive Ballroom",
              "description": "Mobile devices and browsers are now advanced enough that developers can build native-quality mobile apps using open web technologies like HTML5, Javascript, and CSS. In this talk, we’ll provide background on why and how we created Ionic, the design decisions made as we integrated Ionic with Angular, and the performance considerations for mobile platforms that our team had to overcome. We’ll also review new and upcoming Ionic features, and talk about the hidden powers and benefits of combining mobile app development and Angular.",
              "productNames": ["Rachel Rabbit"],
              "timeStart": "9:45 am",
              "timeEnd": "10:00 am",
              "tracks": ["Tooling"],
              "id": "3"
            },
            {
              "name": "University of Ionic",
              "location": "Hall 3",
              "description": "Mobile devices and browsers are now advanced enough that developers can build native-quality mobile apps using open web technologies like HTML5, Javascript, and CSS. In this talk, we’ll provide background on why and how we created Ionic, the design decisions made as we integrated Ionic with Angular, and the performance considerations for mobile platforms that our team had to overcome. We’ll also review new and upcoming Ionic features, and talk about the hidden powers and benefits of combining mobile app development and Angular.",
              "productNames": ["Ellie Elephant"],
              "timeStart": "9:15 am",
              "timeEnd": "9:30 am",
              "tracks": ["Ionic"],
              "id": "4"
            }
          ]
        },
        {
          "time": "10:00 am",
          "offerings": [
            {
              "name": "Coworking startup plan",
              "location": "Hall 1",
              "description": "I want a coworking mobile app that can support #workercount users, in #locationcount place, that can be extended to #extendableusers users in #extendableplacecount places. It should work in #countriescount countries. It should have billing, vendor integration, social interaction facility. It should work in android and ios system",
              "productNames": ["Eva Eagle", "Coworking mobile app"],
              "fields": [
		   {"name":"#workercount", "dispname": "Number of workers", "options": ["10", "50", "100", "200"], "quote": ["100", "200", "100", "80"] },
   {"name":"#locationcount", "dispname": "Number of locations",  "options": ["100", "200"], "quote": []}
			],
              "quoteformula" :  " #workercount * 100 + #locationcount * 1000 ",
              "variablequoteformulas" : [ 
	{"quotename": "simplequote", "quoteformula": "#workercount * 100 + #locationcount * 1000 "},
	{"quotename": "indiaquote", "quoteformula": "#workercount * 200 + #locationcount * 1000 "}],
              "licensehead": "10:00 am",
              "licensebody": "10:00 am",
              "licensebodyvariable": [
	{"licvarname": "maximumlimit", "licdesc": "The user shall not use more than #workercount users and more than #locationcount locations "},
	{"licvarname": "nationlimit", "licdesc": "The user shall use only in nations listed #nationlist "},
	 }],
              "licensetail": "10:00 am",
              "timeStart": "10:00 am",
              "timeEnd": "10:15 am",
              "tracks": ["Ionic"],
              "id": "5"
            },
            {
              "name": "Coworking co-living plan",
              "location": "Hall 1",
              "description": "I want a coworking mobile app that can support 10 users, in 1 place, that can be extended to 100 users in 20 places. It should work in two countries. It should have billing, vendor integration, social interaction facility. It should work in android and ios system",
              "productNames": ["Eva Eagle", "Coworking mobile app"],
              "timeStart": "10:00 am",
              "timeEnd": "10:15 am",
              "tracks": ["Ionic"],
              "id": "19"
            },
            {
              "name": "What's New in Angular",
              "location": "Hall 3",
              "description": "Mobile devices and browsers are now advanced enough that developers can build native-quality mobile apps using open web technologies like HTML5, Javascript, and CSS. In this talk, we’ll provide background on why and how we created Ionic, the design decisions made as we integrated Ionic with Angular, and the performance considerations for mobile platforms that our team had to overcome. We’ll also review new and upcoming Ionic features, and talk about the hidden powers and benefits of combining mobile app development and Angular.",
              "productNames": ["Rachel Rabbit"],
              "timeStart": "10:15 am",
              "timeEnd": "10:30 am",
              "tracks": ["Angular"],
              "id": "6"
            },
            {
              "name": "The Evolution of Ionicons",
              "location": "Hall 2",
              "description": "Mobile devices and browsers are now advanced enough that developers can build native-quality mobile apps using open web technologies like HTML5, Javascript, and CSS. In this talk, we’ll provide background on why and how we created Ionic, the design decisions made as we integrated Ionic with Angular, and the performance considerations for mobile platforms that our team had to overcome. We’ll also review new and upcoming Ionic features, and talk about the hidden powers and benefits of combining mobile app development and Angular.",
              "productNames": ["Isabella Iguana", "Eva Eagle"],
              "timeStart": "10:15 am",
              "timeEnd": "10:30 am",
              "tracks": ["Design"],
              "id": "7"
            },
            {
              "name": "Ionic Pro",
              "location": "Grand Ballroom A",
              "description": "Mobile devices and browsers are now advanced enough that developers can build native-quality mobile apps using open web technologies like HTML5, Javascript, and CSS. In this talk, we’ll provide background on why and how we created Ionic, the design decisions made as we integrated Ionic with Angular, and the performance considerations for mobile platforms that our team had to overcome. We’ll also review new and upcoming Ionic features, and talk about the hidden powers and benefits of combining mobile app development and Angular.",
              "productNames": ["Charlie Cheetah"],
              "timeStart": "10:45 am",
              "timeEnd": "11:00 am",
              "tracks": ["Services"],
              "id": "8"
            }
          ]
        },
        {
          "time": "11:00 am",
          "offerings": [
            {
              "name": "Ionic Workshop",
              "location": "Hall 1",
              "description": "Mobile devices and browsers are now advanced enough that developers can build native-quality mobile apps using open web technologies like HTML5, Javascript, and CSS. In this talk, we’ll provide background on why and how we created Ionic, the design decisions made as we integrated Ionic with Angular, and the performance considerations for mobile platforms that our team had to overcome. We’ll also review new and upcoming Ionic features, and talk about the hidden powers and benefits of combining mobile app development and Angular.",
              "productNames": ["Karl Kitten", "Lionel Lion"],
              "timeStart": "11:00 am",
              "timeEnd": "11:45 am",
              "tracks": ["Workshop"],
              "id": "9"
            },
            {
              "name": "Community Interaction",
              "location": "Hall 3",
              "description": "Mobile devices and browsers are now advanced enough that developers can build native-quality mobile apps using open web technologies like HTML5, Javascript, and CSS. In this talk, we’ll provide background on why and how we created Ionic, the design decisions made as we integrated Ionic with Angular, and the performance considerations for mobile platforms that our team had to overcome. We’ll also review new and upcoming Ionic features, and talk about the hidden powers and benefits of combining mobile app development and Angular.",
              "productNames": ["Lionel Lion", "Gino Giraffe"],
              "timeStart": "11:30 am",
              "timeEnd": "11:50 am",
              "tracks": ["Communication"],
              "id": "10"
            },
            {
              "name": "Navigation in Ionic",
              "location": "Grand Ballroom A",
              "description": "Mobile devices and browsers are now advanced enough that developers can build native-quality mobile apps using open web technologies like HTML5, Javascript, and CSS. In this talk, we’ll provide background on why and how we created Ionic, the design decisions made as we integrated Ionic with Angular, and the performance considerations for mobile platforms that our team had to overcome. We’ll also review new and upcoming Ionic features, and talk about the hidden powers and benefits of combining mobile app development and Angular.",
              "productNames": ["Rachel Rabbit", "Eva Eagle"],
              "timeStart": "11:30 am",
              "timeEnd": "12:00 pm",
              "tracks": ["Navigation"],
              "id": "11"
            }
          ]
        },
        {
          "time": "12:00 pm",
          "offerings": [
            {
              "name": "Lunch",
              "location": "Dining Hall",
              "description": "Come grab lunch with all the Ionic fanatics and talk all things Ionic",
              "timeStart": "12:00 pm",
              "timeEnd": "1:00 pm",
              "tracks": ["Food"],
              "id": "12"
            }
          ]
        },
        {
          "time": "1:00 pm",
          "offerings": [
            {
              "name": "Ionic in the Enterprise",
              "location": "Hall 1",
              "description": "Mobile devices and browsers are now advanced enough that developers can build native-quality mobile apps using open web technologies like HTML5, Javascript, and CSS. In this talk, we’ll provide background on why and how we created Ionic, the design decisions made as we integrated Ionic with Angular, and the performance considerations for mobile platforms that our team had to overcome. We’ll also review new and upcoming Ionic features, and talk about the hidden powers and benefits of combining mobile app development and Angular.",
              "productNames": ["Paul Puppy"],
              "timeStart": "1:00 pm",
              "timeEnd": "1:15 pm",
              "tracks": ["Communication"],
              "id": "13"
            },
            {
              "name": "Ionic Worldwide",
              "location": "Hall 1",
              "description": "Mobile devices and browsers are now advanced enough that developers can build native-quality mobile apps using open web technologies like HTML5, Javascript, and CSS. In this talk, we’ll provide background on why and how we created Ionic, the design decisions made as we integrated Ionic with Angular, and the performance considerations for mobile platforms that our team had to overcome. We’ll also review new and upcoming Ionic features, and talk about the hidden powers and benefits of combining mobile app development and Angular.",
              "productNames": ["Gino Giraffe"],
              "timeStart": "1:15 pm",
              "timeEnd": "1:30 pm",
              "tracks": ["Communication"],
              "id": "14"
            },
            {
              "name": "The Ionic Package",
              "location": "Grand Ballroom B",
              "description": "Mobile devices and browsers are now advanced enough that developers can build native-quality mobile apps using open web technologies like HTML5, Javascript, and CSS. In this talk, we’ll provide background on why and how we created Ionic, the design decisions made as we integrated Ionic with Angular, and the performance considerations for mobile platforms that our team had to overcome. We’ll also review new and upcoming Ionic features, and talk about the hidden powers and benefits of combining mobile app development and Angular.",
              "productNames": ["Molly Mouse", "Burt Bear"],
              "timeStart": "1:30 pm",
              "timeEnd": "2:00 pm",
              "tracks": ["Services"],
              "id": "15"
            }
          ]
        },
        {
          "time": "2:00 pm",
          "offerings": [
            {
              "name": "Push Notifications in Ionic",
              "location": "Hall 2",
              "description": "Mobile devices and browsers are now advanced enough that developers can build native-quality mobile apps using open web technologies like HTML5, Javascript, and CSS. In this talk, we’ll provide background on why and how we created Ionic, the design decisions made as we integrated Ionic with Angular, and the performance considerations for mobile platforms that our team had to overcome. We’ll also review new and upcoming Ionic features, and talk about the hidden powers and benefits of combining mobile app development and Angular.",
              "productNames": ["Burt Bear", "Charlie Cheetah"],
              "timeStart": "2:00 pm",
              "timeEnd": "2:30 pm",
              "tracks": ["Services"],
              "id": "16"
            },
            {
              "name": "Ionic Documentation",
              "location": "Grand Ballroom B",
              "description": "Mobile devices and browsers are now advanced enough that developers can build native-quality mobile apps using open web technologies like HTML5, Javascript, and CSS. In this talk, we’ll provide background on why and how we created Ionic, the design decisions made as we integrated Ionic with Angular, and the performance considerations for mobile platforms that our team had to overcome. We’ll also review new and upcoming Ionic features, and talk about the hidden powers and benefits of combining mobile app development and Angular.",
              "productNames": ["Donald Duck"],
              "timeStart": "2:30 pm",
              "timeEnd": "2:45 pm",
              "tracks": ["Documentation"],
              "id": "17"
            },
            {
              "name": "UX in Ionic",
              "location": "Hall 3",
              "description": "Mobile devices and browsers are now advanced enough that developers can build native-quality mobile apps using open web technologies like HTML5, Javascript, and CSS. In this talk, we’ll provide background on why and how we created Ionic, the design decisions made as we integrated Ionic with Angular, and the performance considerations for mobile platforms that our team had to overcome. We’ll also review new and upcoming Ionic features, and talk about the hidden powers and benefits of combining mobile app development and Angular.",
              "productNames": ["Isabella Iguana", "Ellie Elephant"],
              "timeStart": "2:45 pm",
              "timeEnd": "3:00 pm",
              "tracks": ["Design"],
              "id": "18"
            }
          ]
        },
        {
          "time": "3:00",
          "offerings": [
            {
              "name": "Angular Directives in Ionic",
              "location": "Hall 1",
              "description": "Mobile devices and browsers are now advanced enough that developers can build native-quality mobile apps using open web technologies like HTML5, Javascript, and CSS. In this talk, we’ll provide background on why and how we created Ionic, the design decisions made as we integrated Ionic with Angular, and the performance considerations for mobile platforms that our team had to overcome. We’ll also review new and upcoming Ionic features, and talk about the hidden powers and benefits of combining mobile app development and Angular.",
              "productNames": ["Ted Turtle"],
              "timeStart": "3:00 pm",
              "timeEnd": "3:30 pm",
              "tracks": ["Angular"],
              "id": "19"
            },
            {
              "name": "Mobile States",
              "location": "Hall 2",
              "description": "Mobile devices and browsers are now advanced enough that developers can build native-quality mobile apps using open web technologies like HTML5, Javascript, and CSS. In this talk, we’ll provide background on why and how we created Ionic, the design decisions made as we integrated Ionic with Angular, and the performance considerations for mobile platforms that our team had to overcome. We’ll also review new and upcoming Ionic features, and talk about the hidden powers and benefits of combining mobile app development and Angular.",
              "productNames": ["Rachel Rabbit"],
              "timeStart": "3:30 pm",
              "timeEnd": "3:45 pm",
              "tracks": ["Navigation"],
              "id": "20"
            }
          ]
        }
      ]
    }
  ],

  "products": [
    {
      "name": "Coworking mobile app",
      "profilePic": "/assets/img/products/bear.jpg",
      "twitter": "ionicframework",
      "about": "Burt is a Bear.",
      "location": "Everywhere",
      "email": "burt@example.com",
      "phone": "+1-541-754-3010",
      "id": "1"
    },
    {
      "name": "Coworking space management system ",
      "profilePic": "/assets/img/products/cheetah.jpg",
      "twitter": "ionicframework",
      "about": "Charlie is a Cheetah.",
      "location": "Everywhere",
      "email": "charlie@example.com",
      "phone": "+1-541-754-3010",
      "id": "2"
    },
    {
      "name": "Coworking admin system ",
      "profilePic": "/assets/img/products/duck.jpg",
      "twitter": "ionicframework",
      "about": "Donald is a Duck.",
      "location": "Everywhere",
      "email": "donald@example.com",
      "phone": "+1-541-754-3010",
      "id": "3"
    },
    {
      "name": "Coworking api integration ",
      "profilePic": "/assets/img/products/eagle.jpg",
      "twitter": "ionicframework",
      "about": "Eva is an Eagle.",
      "location": "Everywhere",
      "email": "eva@example.com",
      "phone": "+1-541-754-3010",
      "id": "4"
    },
    {
      "name": "Karl Kitten",
      "profilePic": "/assets/img/products/kitten.jpg",
      "twitter": "ionicframework",
      "about": "Karl is a Kitten.",
      "location": "Everywhere",
      "email": "karl@example.com",
      "phone": "+1-541-754-3010",
      "id": "8"
    },
    {
      "name": "Lionel Lion",
      "profilePic": "/assets/img/products/lion.jpg",
      "twitter": "ionicframework",
      "about": "Lionel is a Lion.",
      "location": "Everywhere",
      "email": "lionel@example.com",
      "phone": "+1-541-754-3010",
      "id": "9"
    },
    {
      "name": "Molly Mouse",
      "profilePic": "/assets/img/products/mouse.jpg",
      "twitter": "ionicframework",
      "about": "Molly is a Mouse.",
      "location": "Everywhere",
      "email": "molly@example.com",
      "phone": "+1-541-754-3010",
      "id": "10"
    },
    {
      "name": "Paul Puppy",
      "profilePic": "/assets/img/products/puppy.jpg",
      "twitter": "ionicframework",
      "about": "Paul is a Puppy.",
      "location": "Everywhere",
      "email": "paul@example.com",
      "phone": "+1-541-754-3010",
      "id": "11"
    },
    {
      "name": "Rachel Rabbit",
      "profilePic": "/assets/img/products/rabbit.jpg",
      "twitter": "ionicframework",
      "about": "Rachel is a Rabbit.",
      "location": "Everywhere",
      "email": "rachel@example.com",
      "phone": "+1-541-754-3010",
      "id": "12"
    },
    {
      "name": "Ted Turtle",
      "profilePic": "/assets/img/products/turtle.jpg",
      "twitter": "ionicframework",
      "about": "Ted is a Turtle.",
      "location": "Everywhere",
      "email": "ted@example.com",
      "phone": "+1-541-754-3010",
      "id": "13"
    }
  ],

  "map": [
    {
      "name": "Monona Terrace Convention Center",
      "lat": 43.071584,
      "lng": -89.38012,
      "center": true
    },
    {
      "name": "Ionic HQ",
      "lat": 43.074395,
      "lng": -89.381056
    },
    {
      "name": "Afterparty - Brocach Irish Pub",
      "lat": 43.07336,
      "lng": -89.38335
    }
  ]
}
